module FlushUnit (
    input  wire  Branch,
    input  wire  Zero,
    output reg   flush
);
endmodule
