module InstructionMemory (
    input  wire [31:0] address,
    output wire [31:0] instruction
);
endmodule
